module program_reg (
  input  wire        clk,
  input  wire        rst_n,
  input  wire        read,
  input  wire        write,
  input  wire [ 7:0] index,
  input  wire [ 7:0] length,
  input  wire [31:0] data,
  output reg  [31:0] order,
  output reg  [ 7:0] len
);

  reg [31:0] record[0:127];

  always @(posedge clk) begin
    if (!rst_n) len <= 0;
    else if (write) len <= length;
    else len <= len;
  end

  always @(posedge clk) begin
    if (!rst_n) order <= 0;
    else begin
      if (read && !write) begin
        if (index > len) order <= 0;
        else begin
          case (index)
            8'd0:    order <= record[0];
            8'd1:    order <= record[1];
            8'd2:    order <= record[2];
            8'd3:    order <= record[3];
            8'd4:    order <= record[4];
            8'd5:    order <= record[5];
            8'd6:    order <= record[6];
            8'd7:    order <= record[7];
            8'd8:    order <= record[8];
            8'd9:    order <= record[9];
            8'd10:   order <= record[10];
            8'd11:   order <= record[11];
            8'd12:   order <= record[12];
            8'd13:   order <= record[13];
            8'd14:   order <= record[14];
            8'd15:   order <= record[15];
            8'd16:   order <= record[16];
            8'd17:   order <= record[17];
            8'd18:   order <= record[18];
            8'd19:   order <= record[19];
            8'd20:   order <= record[20];
            8'd21:   order <= record[21];
            8'd22:   order <= record[22];
            8'd23:   order <= record[23];
            8'd24:   order <= record[24];
            8'd25:   order <= record[25];
            8'd26:   order <= record[26];
            8'd27:   order <= record[27];
            8'd28:   order <= record[28];
            8'd29:   order <= record[29];
            8'd30:   order <= record[30];
            8'd31:   order <= record[31];
            8'd32:   order <= record[32];
            8'd33:   order <= record[33];
            8'd34:   order <= record[34];
            8'd35:   order <= record[35];
            8'd36:   order <= record[36];
            8'd37:   order <= record[37];
            8'd38:   order <= record[38];
            8'd39:   order <= record[39];
            8'd40:   order <= record[40];
            8'd41:   order <= record[41];
            8'd42:   order <= record[42];
            8'd43:   order <= record[43];
            8'd44:   order <= record[44];
            8'd45:   order <= record[45];
            8'd46:   order <= record[46];
            8'd47:   order <= record[47];
            8'd48:   order <= record[48];
            8'd49:   order <= record[49];
            8'd50:   order <= record[50];
            8'd51:   order <= record[51];
            8'd52:   order <= record[52];
            8'd53:   order <= record[53];
            8'd54:   order <= record[54];
            8'd55:   order <= record[55];
            8'd56:   order <= record[56];
            8'd57:   order <= record[57];
            8'd58:   order <= record[58];
            8'd59:   order <= record[59];
            8'd60:   order <= record[60];
            8'd61:   order <= record[61];
            8'd62:   order <= record[62];
            8'd63:   order <= record[63];
            8'd64:   order <= record[64];
            8'd65:   order <= record[65];
            8'd66:   order <= record[66];
            8'd67:   order <= record[67];
            8'd68:   order <= record[68];
            8'd69:   order <= record[69];
            8'd70:   order <= record[70];
            8'd71:   order <= record[71];
            8'd72:   order <= record[72];
            8'd73:   order <= record[73];
            8'd74:   order <= record[74];
            8'd75:   order <= record[75];
            8'd76:   order <= record[76];
            8'd77:   order <= record[77];
            8'd78:   order <= record[78];
            8'd79:   order <= record[79];
            8'd80:   order <= record[80];
            8'd81:   order <= record[81];
            8'd82:   order <= record[82];
            8'd83:   order <= record[83];
            8'd84:   order <= record[84];
            8'd85:   order <= record[85];
            8'd86:   order <= record[86];
            8'd87:   order <= record[87];
            8'd88:   order <= record[88];
            8'd89:   order <= record[89];
            8'd90:   order <= record[90];
            8'd91:   order <= record[91];
            8'd92:   order <= record[92];
            8'd93:   order <= record[93];
            8'd94:   order <= record[94];
            8'd95:   order <= record[95];
            8'd96:   order <= record[96];
            8'd97:   order <= record[97];
            8'd98:   order <= record[98];
            8'd99:   order <= record[99];
            8'd100:  order <= record[100];
            8'd101:  order <= record[101];
            8'd102:  order <= record[102];
            8'd103:  order <= record[103];
            8'd104:  order <= record[104];
            8'd105:  order <= record[105];
            8'd106:  order <= record[106];
            8'd107:  order <= record[107];
            8'd108:  order <= record[108];
            8'd109:  order <= record[109];
            8'd110:  order <= record[110];
            8'd111:  order <= record[111];
            8'd112:  order <= record[112];
            8'd113:  order <= record[113];
            8'd114:  order <= record[114];
            8'd115:  order <= record[115];
            8'd116:  order <= record[116];
            8'd117:  order <= record[117];
            8'd118:  order <= record[118];
            8'd119:  order <= record[119];
            8'd120:  order <= record[120];
            8'd121:  order <= record[121];
            8'd122:  order <= record[122];
            8'd123:  order <= record[123];
            8'd124:  order <= record[124];
            8'd125:  order <= record[125];
            8'd126:  order <= record[126];
            8'd127:  order <= record[127];
            default: order <= 0;
          endcase
        end
      end else order <= 0;
    end
  end

  always @(posedge clk) begin
    if (!rst_n) begin
      record[0]   <= 0;
      record[1]   <= 0;
      record[2]   <= 0;
      record[3]   <= 0;
      record[4]   <= 0;
      record[5]   <= 0;
      record[6]   <= 0;
      record[7]   <= 0;
      record[8]   <= 0;
      record[9]   <= 0;
      record[10]  <= 0;
      record[11]  <= 0;
      record[12]  <= 0;
      record[13]  <= 0;
      record[14]  <= 0;
      record[15]  <= 0;
      record[16]  <= 0;
      record[17]  <= 0;
      record[18]  <= 0;
      record[19]  <= 0;
      record[20]  <= 0;
      record[21]  <= 0;
      record[22]  <= 0;
      record[23]  <= 0;
      record[24]  <= 0;
      record[25]  <= 0;
      record[26]  <= 0;
      record[27]  <= 0;
      record[28]  <= 0;
      record[29]  <= 0;
      record[30]  <= 0;
      record[31]  <= 0;
      record[32]  <= 0;
      record[33]  <= 0;
      record[34]  <= 0;
      record[35]  <= 0;
      record[36]  <= 0;
      record[37]  <= 0;
      record[38]  <= 0;
      record[39]  <= 0;
      record[40]  <= 0;
      record[41]  <= 0;
      record[42]  <= 0;
      record[43]  <= 0;
      record[44]  <= 0;
      record[45]  <= 0;
      record[46]  <= 0;
      record[47]  <= 0;
      record[48]  <= 0;
      record[49]  <= 0;
      record[50]  <= 0;
      record[51]  <= 0;
      record[52]  <= 0;
      record[53]  <= 0;
      record[54]  <= 0;
      record[55]  <= 0;
      record[56]  <= 0;
      record[57]  <= 0;
      record[58]  <= 0;
      record[59]  <= 0;
      record[60]  <= 0;
      record[61]  <= 0;
      record[62]  <= 0;
      record[63]  <= 0;
      record[64]  <= 0;
      record[65]  <= 0;
      record[66]  <= 0;
      record[67]  <= 0;
      record[68]  <= 0;
      record[69]  <= 0;
      record[70]  <= 0;
      record[71]  <= 0;
      record[72]  <= 0;
      record[73]  <= 0;
      record[74]  <= 0;
      record[75]  <= 0;
      record[76]  <= 0;
      record[77]  <= 0;
      record[78]  <= 0;
      record[79]  <= 0;
      record[80]  <= 0;
      record[81]  <= 0;
      record[82]  <= 0;
      record[83]  <= 0;
      record[84]  <= 0;
      record[85]  <= 0;
      record[86]  <= 0;
      record[87]  <= 0;
      record[88]  <= 0;
      record[89]  <= 0;
      record[90]  <= 0;
      record[91]  <= 0;
      record[92]  <= 0;
      record[93]  <= 0;
      record[94]  <= 0;
      record[95]  <= 0;
      record[96]  <= 0;
      record[97]  <= 0;
      record[98]  <= 0;
      record[99]  <= 0;
      record[100] <= 0;
      record[101] <= 0;
      record[102] <= 0;
      record[103] <= 0;
      record[104] <= 0;
      record[105] <= 0;
      record[106] <= 0;
      record[107] <= 0;
      record[108] <= 0;
      record[109] <= 0;
      record[110] <= 0;
      record[111] <= 0;
      record[112] <= 0;
      record[113] <= 0;
      record[114] <= 0;
      record[115] <= 0;
      record[116] <= 0;
      record[117] <= 0;
      record[118] <= 0;
      record[119] <= 0;
      record[120] <= 0;
      record[121] <= 0;
      record[122] <= 0;
      record[123] <= 0;
      record[124] <= 0;
      record[125] <= 0;
      record[126] <= 0;
      record[127] <= 0;
    end else begin
      if (!write) begin
        record[0]   <= record[0];
        record[1]   <= record[1];
        record[2]   <= record[2];
        record[3]   <= record[3];
        record[4]   <= record[4];
        record[5]   <= record[5];
        record[6]   <= record[6];
        record[7]   <= record[7];
        record[8]   <= record[8];
        record[9]   <= record[9];
        record[10]  <= record[10];
        record[11]  <= record[11];
        record[12]  <= record[12];
        record[13]  <= record[13];
        record[14]  <= record[14];
        record[15]  <= record[15];
        record[16]  <= record[16];
        record[17]  <= record[17];
        record[18]  <= record[18];
        record[19]  <= record[19];
        record[20]  <= record[20];
        record[21]  <= record[21];
        record[22]  <= record[22];
        record[23]  <= record[23];
        record[24]  <= record[24];
        record[25]  <= record[25];
        record[26]  <= record[26];
        record[27]  <= record[27];
        record[28]  <= record[28];
        record[29]  <= record[29];
        record[30]  <= record[30];
        record[31]  <= record[31];
        record[32]  <= record[32];
        record[33]  <= record[33];
        record[34]  <= record[34];
        record[35]  <= record[35];
        record[36]  <= record[36];
        record[37]  <= record[37];
        record[38]  <= record[38];
        record[39]  <= record[39];
        record[40]  <= record[40];
        record[41]  <= record[41];
        record[42]  <= record[42];
        record[43]  <= record[43];
        record[44]  <= record[44];
        record[45]  <= record[45];
        record[46]  <= record[46];
        record[47]  <= record[47];
        record[48]  <= record[48];
        record[49]  <= record[49];
        record[50]  <= record[50];
        record[51]  <= record[51];
        record[52]  <= record[52];
        record[53]  <= record[53];
        record[54]  <= record[54];
        record[55]  <= record[55];
        record[56]  <= record[56];
        record[57]  <= record[57];
        record[58]  <= record[58];
        record[59]  <= record[59];
        record[60]  <= record[60];
        record[61]  <= record[61];
        record[62]  <= record[62];
        record[63]  <= record[63];
        record[64]  <= record[64];
        record[65]  <= record[65];
        record[66]  <= record[66];
        record[67]  <= record[67];
        record[68]  <= record[68];
        record[69]  <= record[69];
        record[70]  <= record[70];
        record[71]  <= record[71];
        record[72]  <= record[72];
        record[73]  <= record[73];
        record[74]  <= record[74];
        record[75]  <= record[75];
        record[76]  <= record[76];
        record[77]  <= record[77];
        record[78]  <= record[78];
        record[79]  <= record[79];
        record[80]  <= record[80];
        record[81]  <= record[81];
        record[82]  <= record[82];
        record[83]  <= record[83];
        record[84]  <= record[84];
        record[85]  <= record[85];
        record[86]  <= record[86];
        record[87]  <= record[87];
        record[88]  <= record[88];
        record[89]  <= record[89];
        record[90]  <= record[90];
        record[91]  <= record[91];
        record[92]  <= record[92];
        record[93]  <= record[93];
        record[94]  <= record[94];
        record[95]  <= record[95];
        record[96]  <= record[96];
        record[97]  <= record[97];
        record[98]  <= record[98];
        record[99]  <= record[99];
        record[100] <= record[100];
        record[101] <= record[101];
        record[102] <= record[102];
        record[103] <= record[103];
        record[104] <= record[104];
        record[105] <= record[105];
        record[106] <= record[106];
        record[107] <= record[107];
        record[108] <= record[108];
        record[109] <= record[109];
        record[110] <= record[110];
        record[111] <= record[111];
        record[112] <= record[112];
        record[113] <= record[113];
        record[114] <= record[114];
        record[115] <= record[115];
        record[116] <= record[116];
        record[117] <= record[117];
        record[118] <= record[118];
        record[119] <= record[119];
        record[120] <= record[120];
        record[121] <= record[121];
        record[122] <= record[122];
        record[123] <= record[123];
        record[124] <= record[124];
        record[125] <= record[125];
        record[126] <= record[126];
        record[127] <= record[127];
      end else
        case (index)
          8'd0:   record[0] <= data;
          8'd1:   record[1] <= data;
          8'd2:   record[2] <= data;
          8'd3:   record[3] <= data;
          8'd4:   record[4] <= data;
          8'd5:   record[5] <= data;
          8'd6:   record[6] <= data;
          8'd7:   record[7] <= data;
          8'd8:   record[8] <= data;
          8'd9:   record[9] <= data;
          8'd10:  record[10] <= data;
          8'd11:  record[11] <= data;
          8'd12:  record[12] <= data;
          8'd13:  record[13] <= data;
          8'd14:  record[14] <= data;
          8'd15:  record[15] <= data;
          8'd16:  record[16] <= data;
          8'd17:  record[17] <= data;
          8'd18:  record[18] <= data;
          8'd19:  record[19] <= data;
          8'd20:  record[20] <= data;
          8'd21:  record[21] <= data;
          8'd22:  record[22] <= data;
          8'd23:  record[23] <= data;
          8'd24:  record[24] <= data;
          8'd25:  record[25] <= data;
          8'd26:  record[26] <= data;
          8'd27:  record[27] <= data;
          8'd28:  record[28] <= data;
          8'd29:  record[29] <= data;
          8'd30:  record[30] <= data;
          8'd31:  record[31] <= data;
          8'd32:  record[32] <= data;
          8'd33:  record[33] <= data;
          8'd34:  record[34] <= data;
          8'd35:  record[35] <= data;
          8'd36:  record[36] <= data;
          8'd37:  record[37] <= data;
          8'd38:  record[38] <= data;
          8'd39:  record[39] <= data;
          8'd40:  record[40] <= data;
          8'd41:  record[41] <= data;
          8'd42:  record[42] <= data;
          8'd43:  record[43] <= data;
          8'd44:  record[44] <= data;
          8'd45:  record[45] <= data;
          8'd46:  record[46] <= data;
          8'd47:  record[47] <= data;
          8'd48:  record[48] <= data;
          8'd49:  record[49] <= data;
          8'd50:  record[50] <= data;
          8'd51:  record[51] <= data;
          8'd52:  record[52] <= data;
          8'd53:  record[53] <= data;
          8'd54:  record[54] <= data;
          8'd55:  record[55] <= data;
          8'd56:  record[56] <= data;
          8'd57:  record[57] <= data;
          8'd58:  record[58] <= data;
          8'd59:  record[59] <= data;
          8'd60:  record[60] <= data;
          8'd61:  record[61] <= data;
          8'd62:  record[62] <= data;
          8'd63:  record[63] <= data;
          8'd64:  record[64] <= data;
          8'd65:  record[65] <= data;
          8'd66:  record[66] <= data;
          8'd67:  record[67] <= data;
          8'd68:  record[68] <= data;
          8'd69:  record[69] <= data;
          8'd70:  record[70] <= data;
          8'd71:  record[71] <= data;
          8'd72:  record[72] <= data;
          8'd73:  record[73] <= data;
          8'd74:  record[74] <= data;
          8'd75:  record[75] <= data;
          8'd76:  record[76] <= data;
          8'd77:  record[77] <= data;
          8'd78:  record[78] <= data;
          8'd79:  record[79] <= data;
          8'd80:  record[80] <= data;
          8'd81:  record[81] <= data;
          8'd82:  record[82] <= data;
          8'd83:  record[83] <= data;
          8'd84:  record[84] <= data;
          8'd85:  record[85] <= data;
          8'd86:  record[86] <= data;
          8'd87:  record[87] <= data;
          8'd88:  record[88] <= data;
          8'd89:  record[89] <= data;
          8'd90:  record[90] <= data;
          8'd91:  record[91] <= data;
          8'd92:  record[92] <= data;
          8'd93:  record[93] <= data;
          8'd94:  record[94] <= data;
          8'd95:  record[95] <= data;
          8'd96:  record[96] <= data;
          8'd97:  record[97] <= data;
          8'd98:  record[98] <= data;
          8'd99:  record[99] <= data;
          8'd100: record[100] <= data;
          8'd101: record[101] <= data;
          8'd102: record[102] <= data;
          8'd103: record[103] <= data;
          8'd104: record[104] <= data;
          8'd105: record[105] <= data;
          8'd106: record[106] <= data;
          8'd107: record[107] <= data;
          8'd108: record[108] <= data;
          8'd109: record[109] <= data;
          8'd110: record[110] <= data;
          8'd111: record[111] <= data;
          8'd112: record[112] <= data;
          8'd113: record[113] <= data;
          8'd114: record[114] <= data;
          8'd115: record[115] <= data;
          8'd116: record[116] <= data;
          8'd117: record[117] <= data;
          8'd118: record[118] <= data;
          8'd119: record[119] <= data;
          8'd120: record[120] <= data;
          8'd121: record[121] <= data;
          8'd122: record[122] <= data;
          8'd123: record[123] <= data;
          8'd124: record[124] <= data;
          8'd125: record[125] <= data;
          8'd126: record[126] <= data;
          8'd127: record[127] <= data;
          default: begin
            record[0]   <= record[0];
            record[1]   <= record[1];
            record[2]   <= record[2];
            record[3]   <= record[3];
            record[4]   <= record[4];
            record[5]   <= record[5];
            record[6]   <= record[6];
            record[7]   <= record[7];
            record[8]   <= record[8];
            record[9]   <= record[9];
            record[10]  <= record[10];
            record[11]  <= record[11];
            record[12]  <= record[12];
            record[13]  <= record[13];
            record[14]  <= record[14];
            record[15]  <= record[15];
            record[16]  <= record[16];
            record[17]  <= record[17];
            record[18]  <= record[18];
            record[19]  <= record[19];
            record[20]  <= record[20];
            record[21]  <= record[21];
            record[22]  <= record[22];
            record[23]  <= record[23];
            record[24]  <= record[24];
            record[25]  <= record[25];
            record[26]  <= record[26];
            record[27]  <= record[27];
            record[28]  <= record[28];
            record[29]  <= record[29];
            record[30]  <= record[30];
            record[31]  <= record[31];
            record[32]  <= record[32];
            record[33]  <= record[33];
            record[34]  <= record[34];
            record[35]  <= record[35];
            record[36]  <= record[36];
            record[37]  <= record[37];
            record[38]  <= record[38];
            record[39]  <= record[39];
            record[40]  <= record[40];
            record[41]  <= record[41];
            record[42]  <= record[42];
            record[43]  <= record[43];
            record[44]  <= record[44];
            record[45]  <= record[45];
            record[46]  <= record[46];
            record[47]  <= record[47];
            record[48]  <= record[48];
            record[49]  <= record[49];
            record[50]  <= record[50];
            record[51]  <= record[51];
            record[52]  <= record[52];
            record[53]  <= record[53];
            record[54]  <= record[54];
            record[55]  <= record[55];
            record[56]  <= record[56];
            record[57]  <= record[57];
            record[58]  <= record[58];
            record[59]  <= record[59];
            record[60]  <= record[60];
            record[61]  <= record[61];
            record[62]  <= record[62];
            record[63]  <= record[63];
            record[64]  <= record[64];
            record[65]  <= record[65];
            record[66]  <= record[66];
            record[67]  <= record[67];
            record[68]  <= record[68];
            record[69]  <= record[69];
            record[70]  <= record[70];
            record[71]  <= record[71];
            record[72]  <= record[72];
            record[73]  <= record[73];
            record[74]  <= record[74];
            record[75]  <= record[75];
            record[76]  <= record[76];
            record[77]  <= record[77];
            record[78]  <= record[78];
            record[79]  <= record[79];
            record[80]  <= record[80];
            record[81]  <= record[81];
            record[82]  <= record[82];
            record[83]  <= record[83];
            record[84]  <= record[84];
            record[85]  <= record[85];
            record[86]  <= record[86];
            record[87]  <= record[87];
            record[88]  <= record[88];
            record[89]  <= record[89];
            record[90]  <= record[90];
            record[91]  <= record[91];
            record[92]  <= record[92];
            record[93]  <= record[93];
            record[94]  <= record[94];
            record[95]  <= record[95];
            record[96]  <= record[96];
            record[97]  <= record[97];
            record[98]  <= record[98];
            record[99]  <= record[99];
            record[100] <= record[100];
            record[101] <= record[101];
            record[102] <= record[102];
            record[103] <= record[103];
            record[104] <= record[104];
            record[105] <= record[105];
            record[106] <= record[106];
            record[107] <= record[107];
            record[108] <= record[108];
            record[109] <= record[109];
            record[110] <= record[110];
            record[111] <= record[111];
            record[112] <= record[112];
            record[113] <= record[113];
            record[114] <= record[114];
            record[115] <= record[115];
            record[116] <= record[116];
            record[117] <= record[117];
            record[118] <= record[118];
            record[119] <= record[119];
            record[120] <= record[120];
            record[121] <= record[121];
            record[122] <= record[122];
            record[123] <= record[123];
            record[124] <= record[124];
            record[125] <= record[125];
            record[126] <= record[126];
            record[127] <= record[127];
          end
        endcase
    end
  end

endmodule
