module counter_16bit();
endmodule